.include gpdk90nm_tt.cir

* PARAMS * TODO: change:
.param ln = 350n 
.param lp = 350n
.param wn = 700n
.param wp = 1500n

.param VDD = 1V
.param VSS = 0V



*********************
* TRANSMISSION GATE *
*********************

*       name                input   pmos gate   nmos gate   output  powerup powerdown
.subckt transmission_gate   inp     pmos_gate   nmos_gate   outp    VDD     VSS

*           Drain   Gate        Source  Bulk    Type    Length  Width
internal_p1 outp    pmos_gate   inp     VDD     pmos1v  l = lp  w = wp
internal_n1 inp     nmos_gate   outp    VSS     nmos1v  l = ln  w = wn

.ends



************
* NOT GATE *
************

*       name     input  output  powerup powerdown
.subckt not_gate inp    outp    VDD     VSS

*           Drain   Gate    Source  Bulk    Type   Length   Width
internal_p2 outp    inp     VDD     VDD     pmos1v l = lp   w = wp
internal_n2 outp    inp     VSS     VSS     nmos1v l = ln   w = wn

.ends



***********
* BITCELL *
***********

*       name    input   output  writeEN     writeENneg  readEN      readENneg   powerup powerdown
.subckt bitcell inp     outp    we          wen         re          ren         VDD     VSS

* kanskje TODO: definer Q0, Q1, Q2

*   input   pmos gate   nmos gate   output  powerup powerdown   type(transmission_gate)
TG1 inp     wen         we          Q0      VDD     VSS         transmission_gate
TG2 Q2      we          wen         Q0      VDD     VSS         transmission_gate
TG3 Q2      ren         re          outp    VDD     VSS         transmission_gate

*       input   output  powerup powerdown   type(not_gate)
NOT1    Q0      Q1      VDD     VSS         not_gate
NOT2    Q1      Q2      VDD     VSS         not_gate

.ends



*********
* SIMUL *
*********

*   input   output  writeEN     writeENneg  readEN      readENneg   powerup powerdown   type(bitcell)
BC1 data    outp    we          wen         re          ren         VDD     VSS         bitcell

.dc data 0 1 0.01

